module register_addressing(
  input wire [27:0] instruction,
  output wire [3:0] Rn, Rm, Rs
);

endmodule
